/* Types are defined here for all other Bluespec files to include */

package types;

import MIPS1_Instruction32::*;

`define Instruction_OpCode MIPS1_Instruction_Opcode;

endpackage
